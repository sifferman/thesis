
assign out =
    in[31] ? 31 : in[30] ? 30 :
    in[29] ? 29 : in[28] ? 28 :
    in[27] ? 27 : in[26] ? 26 :
    in[25] ? 25 : in[24] ? 24 :
    in[23] ? 23 : in[22] ? 22 :
    in[21] ? 21 : in[20] ? 20 :
    in[19] ? 19 : in[18] ? 18 :
    in[17] ? 17 : in[16] ? 16 :
    in[15] ? 15 : in[14] ? 14 :
    in[13] ? 13 : in[12] ? 12 :
    in[11] ? 11 : in[10] ? 10 :
    in[ 9] ?  9 : in[ 8] ?  8 :
    in[ 7] ?  7 : in[ 6] ?  6 :
    in[ 5] ?  5 : in[ 4] ?  4 :
    in[ 3] ?  3 : in[ 2] ?  2 :
    in[ 1] ?  1 : 0;
